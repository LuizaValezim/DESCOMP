library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Decoder is
	port (
		OPCODE : in std_logic_vector(5 downto 0);
		FUNCT : in std_logic_vector(5 downto 0);
		OPERACAO : in std_logic_vector(1 downto 0);
		outPUT : out std_logic_vector(8 downto 0)
	);
end entity;

architecture arch_name OF Decoder is
	constant ADDR : std_logic_vector(5 downto 0) := "100000";
	constant SUBR : std_logic_vector(5 downto 0) := "100010";
	constant LW : std_logic_vector(5 downto 0) := "100011";
	constant SW : std_logic_vector(5 downto 0) := "101011";
	constant BEQ : std_logic_vector(5 downto 0) := "000100";
	constant J : std_logic_vector(5 downto 0) := "000010";
	constant SLT : std_logic_vector(5 downto 0) := "101010";
	constant ANDR : std_logic_vector(5 downto 0) := "100100";
	constant ORR : std_logic_vector(5 downto 0) := "100101";

begin

	outPUT <= "0" & "0011"  & "1010" when (OPCODE = LW) else
		"0" & "0001"   & "0001" when (OPCODE = SW) else
		"0" & "0000"  & "0100" when (OPCODE = BEQ) else
		"1" & "0110"  & "0000" when (((FUNCT = ADDR) OR (FUNCT = SUBR) OR (FUNCT = ORR) OR (FUNCT = ANDR) OR (FUNCT = SLT)) AND OPCODE = "000000") else
		"0" & "1000"  & "0000" when (OPCODE = J) else
		"000000000";
end architecture;