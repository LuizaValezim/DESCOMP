library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 15;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (8 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI : std_logic_vector(3 downto 0) := "0100";
  constant STA : std_logic_vector(3 downto 0) := "0101";
  constant JMP : std_logic_vector(3 downto 0) := "0110";
  constant JEQ : std_logic_vector(3 downto 0) := "0111";
  constant CEQ : std_logic_vector(3 downto 0) := "1000";
  constant JSR : std_logic_vector(3 downto 0) := "1001";
  constant RET : std_logic_vector(3 downto 0) := "1010";
  constant ANDI : std_logic_vector(3 downto 0) := "1011";
  constant CLT : std_logic_vector (3 downto 0) := "1100"; 
  constant JLT : std_logic_vector (3 downto 0) := "1101"; 
  constant ADDI : std_logic_vector (3 downto 0) := "1110"; 
  constant R0:    std_logic_vector (1 DOWNTO 0)	:= "00";
  constant R1:    std_logic_vector (1 DOWNTO 0)	:= "01";
  constant R2:    std_logic_vector (1 DOWNTO 0)	:= "10";
  constant R3:    std_logic_vector (1 DOWNTO 0)	:= "11";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
		
  begin
		tmp(0) := LDI  &  R0  &  '0'  &  x"00";	    
		tmp(1) := LDI  &  R1  &  '0'  &  x"01";	    
		tmp(2) := LDI  &  R2  &  '0'  &  x"06";	    
		tmp(3) := LDI  &  R3  &  '0'  &  x"0a";	    
		tmp(7) := STA  &  R0  &  '1'  &  x"20";	    
		tmp(8) := STA  &  R0  &  '1'  &  x"21";	    
		tmp(9) := STA  &  R0  &  '1'  &  x"22";	    
		tmp(10) := STA  &  R0  &  '1'  &  x"23";	
		tmp(11) := STA  &  R0  &  '1'  &  x"24";	
		tmp(12) := STA  &  R0  &  '1'  &  x"25";	
		tmp(13) := STA  &  R0  &  '0'  &  x"00";	
		tmp(14) := STA  &  R0  &  '0'  &  x"01";	
		tmp(15) := STA  &  R0  &  '0'  &  x"02";	
		tmp(16) := STA  &  R0  &  '0'  &  x"03";	
		tmp(17) := STA  &  R0  &  '0'  &  x"04";	
		tmp(18) := STA  &  R0  &  '0'  &  x"05";	
		tmp(20) := STA  &  R0  &  '0'  &  x"07";	
		tmp(21) := STA  &  R1  &  '0'  &  x"08";	
		tmp(22) := STA  &  R3  &  '0'  &  x"09";	
		tmp(29) := STA  &  R2  &  '0'  &  x"10";	
		tmp(30) := LDI  &  R0  &  '0'  &  x"02";	
		tmp(31) := STA  &  R0  &  '0'  &  x"11";	
		tmp(32) := LDI  &  R0  &  '0'  &  x"04";	
		tmp(33) := STA  &  R0  &  '0'  &  x"12";	
		tmp(34) := LDI  &  R0  &  '0'  &  x"18";	
		tmp(35) := STA  &  R0  &  '0'  &  x"13";	
		tmp(36) := NOP  &  R0  &  '0'  &  x"00";	
		tmp(37) := LDA  &  R0  &  '1'  &  x"60";	
		tmp(38) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(39) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(40) := JEQ  &  R0  &  '0'  &  x"2b";	
		tmp(41) := JSR  &  R0  &  '0'  &  x"45";	
		tmp(42) := NOP  &  R0  &  '0'  &  x"00";	
		tmp(43) := LDA  &  R1  &  '1'  &  x"61";	
		tmp(44) := ANDI  &  R1  &  '0'  &  x"01";	
		tmp(45) := CEQ  &  R1  &  '0'  &  x"07";	
		tmp(46) := JEQ  &  R0  &  '0'  &  x"31";	
		tmp(47) := JSR  &  R0  &  '0'  &  x"bb";	
		tmp(48) := NOP  &  R0  &  '0'  &  x"00";	
		tmp(49) := JSR  &  R0  &  '0'  &  x"a0";	
		tmp(50) := NOP  &  R0  &  '0'  &  x"00";	
		tmp(51) := LDA  &  R0  &  '1'  &  x"62";	
		tmp(52) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(53) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(54) := JEQ  &  R0  &  '0'  &  x"38";	
		tmp(55) := JSR  &  R0  &  '1'  &  x"28";	
		tmp(56) := LDA  &  R2  &  '1'  &  x"63";	
		tmp(57) := ANDI  &  R2  &  '0'  &  x"01";	
		tmp(58) := CEQ  &  R2  &  '0'  &  x"07";	
		tmp(59) := JEQ  &  R0  &  '0'  &  x"3e";	
		tmp(60) := JSR  &  R0  &  '1'  &  x"35";	
		tmp(61) := NOP  &  R0  &  '0'  &  x"00";	
		tmp(62) := LDA  &  R3  &  '1'  &  x"64";	
		tmp(63) := ANDI  &  R3  &  '0'  &  x"01";	
		tmp(64) := CEQ  &  R3  &  '0'  &  x"08";	
		tmp(65) := JEQ  &  R0  &  '0'  &  x"43";	
		tmp(66) := JSR  &  R0  &  '0'  &  x"95";	
		tmp(67) := JSR  &  R0  &  '0'  &  x"83";	
		tmp(68) := JMP  &  R0  &  '0'  &  x"24";	
		tmp(69) := STA  &  R0  &  '1'  &  x"ff";	
		tmp(70) := LDA  &  R0  &  '0'  &  x"00";	
		tmp(71) := ADDI  &  R0  &  '0'  &  x"01";	
		tmp(72) := CEQ  &  R0  &  '0'  &  x"09";	
		tmp(73) := JEQ  &  R0  &  '0'  &  x"4c";	
		tmp(74) := STA  &  R0  &  '0'  &  x"00";	
		tmp(75) := JMP  &  R0  &  '0'  &  x"82";	
		tmp(76) := LDA  &  R0  &  '0'  &  x"07";	
		tmp(77) := STA  &  R0  &  '0'  &  x"00";	
		tmp(78) := LDA  &  R0  &  '0'  &  x"01";	
		tmp(79) := ADDI  &  R0  &  '0'  &  x"01";	
		tmp(80) := CEQ  &  R0  &  '0'  &  x"10";	
		tmp(81) := JEQ  &  R0  &  '0'  &  x"54";	
		tmp(82) := STA  &  R0  &  '0'  &  x"01";	
		tmp(83) := JMP  &  R0  &  '0'  &  x"82";	
		tmp(84) := LDA  &  R0  &  '0'  &  x"07";	
		tmp(85) := STA  &  R0  &  '0'  &  x"01";	
		tmp(86) := LDA  &  R0  &  '0'  &  x"02";	
		tmp(87) := ADDI  &  R0  &  '0'  &  x"01";	
		tmp(88) := CEQ  &  R0  &  '0'  &  x"09";	
		tmp(89) := JEQ  &  R0  &  '0'  &  x"5c";	
		tmp(90) := STA  &  R0  &  '0'  &  x"02";	
		tmp(91) := JMP  &  R0  &  '0'  &  x"82";	
		tmp(92) := LDA  &  R0  &  '0'  &  x"07";	
		tmp(93) := STA  &  R0  &  '0'  &  x"02";	
		tmp(94) := LDA  &  R0  &  '0'  &  x"03";	
		tmp(95) := ADDI  &  R0  &  '0'  &  x"01";	
		tmp(96) := CEQ  &  R0  &  '0'  &  x"10";	
		tmp(97) := JEQ  &  R0  &  '0'  &  x"64";	
		tmp(98) := STA  &  R0  &  '0'  &  x"03";	
		tmp(99) := JMP  &  R0  &  '0'  &  x"82";	
		tmp(100) := LDA  &  R0  &  '0'  &  x"07";	
		tmp(101) := STA  &  R0  &  '0'  &  x"03";	
		tmp(102) := LDA  &  R0  &  '0'  &  x"04";	
		tmp(103) := ADDI  &  R0  &  '0'  &  x"01";	
		tmp(104) := CEQ  &  R0  &  '0'  &  x"12";	
		tmp(105) := JEQ  &  R0  &  '0'  &  x"6e";	
		tmp(106) := CEQ  &  R0  &  '0'  &  x"09";	
		tmp(107) := JEQ  &  R0  &  '0'  &  x"75";	
		tmp(108) := STA  &  R0  &  '0'  &  x"04";	
		tmp(109) := JMP  &  R0  &  '0'  &  x"82";	
		tmp(110) := LDA  &  R1  &  '0'  &  x"05";	
		tmp(111) := CEQ  &  R1  &  '0'  &  x"11";	
		tmp(112) := JEQ  &  R0  &  '0'  &  x"7b";	
		tmp(113) := CEQ  &  R0  &  '0'  &  x"09";	
		tmp(114) := JEQ  &  R0  &  '0'  &  x"75";	
		tmp(115) := STA  &  R0  &  '0'  &  x"04";	
		tmp(116) := JMP  &  R0  &  '0'  &  x"82";	
		tmp(117) := LDA  &  R0  &  '0'  &  x"07";	
		tmp(118) := STA  &  R0  &  '0'  &  x"04";	
		tmp(119) := LDA  &  R0  &  '0'  &  x"05";	
		tmp(120) := ADDI  &  R0  &  '0'  &  x"01";	
		tmp(121) := STA  &  R0  &  '0'  &  x"05";	
		tmp(122) := JMP  &  R0  &  '0'  &  x"82";	
		tmp(123) := LDA  &  R0  &  '0'  &  x"07";	
		tmp(124) := STA  &  R0  &  '0'  &  x"00";	
		tmp(125) := STA  &  R0  &  '0'  &  x"01";	
		tmp(126) := STA  &  R0  &  '0'  &  x"02";	
		tmp(127) := STA  &  R0  &  '0'  &  x"03";	
		tmp(128) := STA  &  R0  &  '0'  &  x"04";	
		tmp(129) := STA  &  R0  &  '0'  &  x"05";	
		tmp(130) := RET  &  R0  &  '0'  &  x"00";	
		tmp(131) := LDA  &  R0  &  '0'  &  x"00";	
		tmp(132) := LDA  &  R1  &  '0'  &  x"01";	
		tmp(133) := LDA  &  R2  &  '0'  &  x"02";	
		tmp(134) := STA  &  R0  &  '1'  &  x"20";	
		tmp(135) := STA  &  R1  &  '1'  &  x"21";	
		tmp(136) := STA  &  R2  &  '1'  &  x"22";	
		tmp(137) := LDA  &  R0  &  '0'  &  x"03";	
		tmp(138) := LDA  &  R1  &  '0'  &  x"04";	
		tmp(139) := LDA  &  R2  &  '0'  &  x"05";	
		tmp(140) := STA  &  R0  &  '1'  &  x"23";	
		tmp(141) := STA  &  R1  &  '1'  &  x"24";	
		tmp(142) := STA  &  R2  &  '1'  &  x"25";	
		tmp(143) := LDA  &  R0  &  '0'  &  x"06";	
		tmp(144) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(145) := JEQ  &  R0  &  '0'  &  x"94";	
		tmp(146) := LDA  &  R2  &  '0'  &  x"08";	
		tmp(148) := RET  &  R0  &  '0'  &  x"00";	
		tmp(149) := LDA  &  R0  &  '0'  &  x"07";	
		tmp(150) := STA  &  R0  &  '0'  &  x"00";	
		tmp(151) := STA  &  R0  &  '0'  &  x"01";	
		tmp(152) := STA  &  R0  &  '0'  &  x"02";	
		tmp(153) := STA  &  R0  &  '0'  &  x"03";	
		tmp(154) := STA  &  R0  &  '0'  &  x"04";	
		tmp(155) := STA  &  R0  &  '0'  &  x"05";	
		tmp(159) := RET  &  R0  &  '0'  &  x"00";	
		tmp(160) := LDA  &  R0  &  '0'  &  x"0a";	
		tmp(161) := CEQ  &  R0  &  '0'  &  x"00";	
		tmp(162) := JEQ  &  R0  &  '0'  &  x"a4";	
		tmp(163) := JMP  &  R0  &  '0'  &  x"ba";	
		tmp(164) := LDA  &  R1  &  '0'  &  x"0b";	
		tmp(165) := CEQ  &  R1  &  '0'  &  x"01";	
		tmp(166) := JEQ  &  R0  &  '0'  &  x"a8";	
		tmp(167) := JMP  &  R0  &  '0'  &  x"ba";	
		tmp(168) := LDA  &  R2  &  '0'  &  x"0c";	
		tmp(169) := CEQ  &  R2  &  '0'  &  x"02";	
		tmp(170) := JEQ  &  R0  &  '0'  &  x"ac";	
		tmp(171) := JMP  &  R0  &  '0'  &  x"ba";	
		tmp(172) := LDA  &  R3  &  '0'  &  x"0d";	
		tmp(173) := CEQ  &  R3  &  '0'  &  x"03";	
		tmp(174) := JEQ  &  R0  &  '0'  &  x"b0";	
		tmp(175) := JMP  &  R0  &  '0'  &  x"ba";	
		tmp(176) := LDA  &  R0  &  '0'  &  x"0e";	
		tmp(177) := CEQ  &  R0  &  '0'  &  x"04";	
		tmp(178) := JEQ  &  R0  &  '0'  &  x"b4";	
		tmp(179) := JMP  &  R0  &  '0'  &  x"ba";	
		tmp(180) := LDA  &  R1  &  '0'  &  x"0f";	
		tmp(181) := CEQ  &  R1  &  '0'  &  x"05";	
		tmp(182) := JEQ  &  R0  &  '0'  &  x"b8";	
		tmp(183) := JMP  &  R0  &  '0'  &  x"ba";	
		tmp(184) := LDA  &  R2  &  '0'  &  x"08";	
		tmp(186) := RET  &  R0  &  '0'  &  x"00";	
		tmp(187) := STA  &  R0  &  '1'  &  x"fe";	
		tmp(190) := JEQ  &  R0  &  '0'  &  x"c2";	
		tmp(191) := LDA  &  R3  &  '0'  &  x"07";	
		tmp(194) := LDA  &  R1  &  '0'  &  x"08";	
		tmp(196) := LDA  &  R0  &  '1'  &  x"61";	
		tmp(197) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(198) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(199) := LDA  &  R2  &  '1'  &  x"40";	
		tmp(200) := JEQ  &  R0  &  '0'  &  x"c2";	
		tmp(201) := STA  &  R2  &  '0'  &  x"0a";	
		tmp(202) := STA  &  R2  &  '1'  &  x"20";	
		tmp(203) := STA  &  R0  &  '1'  &  x"fe";	
		tmp(204) := LDI  &  R1  &  '0'  &  x"02";	
		tmp(206) := LDA  &  R0  &  '1'  &  x"61";	
		tmp(207) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(208) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(209) := LDA  &  R2  &  '1'  &  x"40";	
		tmp(210) := JEQ  &  R0  &  '0'  &  x"cc";	
		tmp(211) := STA  &  R2  &  '0'  &  x"0b";	
		tmp(212) := STA  &  R2  &  '1'  &  x"21";	
		tmp(213) := STA  &  R0  &  '1'  &  x"fe";	
		tmp(214) := LDI  &  R1  &  '0'  &  x"04";	
		tmp(216) := LDA  &  R0  &  '1'  &  x"61";	
		tmp(217) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(218) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(219) := LDA  &  R2  &  '1'  &  x"40";	
		tmp(220) := JEQ  &  R0  &  '0'  &  x"d6";	
		tmp(221) := STA  &  R2  &  '0'  &  x"0c";	
		tmp(222) := STA  &  R2  &  '1'  &  x"22";	
		tmp(223) := STA  &  R0  &  '1'  &  x"fe";	
		tmp(224) := LDI  &  R1  &  '0'  &  x"08";	
		tmp(226) := LDA  &  R0  &  '1'  &  x"61";	
		tmp(227) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(228) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(229) := LDA  &  R2  &  '1'  &  x"40";	
		tmp(230) := JEQ  &  R0  &  '0'  &  x"e0";	
		tmp(231) := STA  &  R2  &  '0'  &  x"0d";	
		tmp(232) := STA  &  R2  &  '1'  &  x"23";	
		tmp(233) := STA  &  R0  &  '1'  &  x"fe";	
		tmp(234) := LDI  &  R1  &  '0'  &  x"10";	
		tmp(236) := LDA  &  R0  &  '1'  &  x"61";	
		tmp(237) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(238) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(239) := LDA  &  R2  &  '1'  &  x"40";	
		tmp(240) := JEQ  &  R0  &  '0'  &  x"ea";	
		tmp(241) := STA  &  R2  &  '0'  &  x"0e";	
		tmp(242) := STA  &  R2  &  '1'  &  x"24";	
		tmp(243) := STA  &  R0  &  '1'  &  x"fe";	
		tmp(244) := LDI  &  R1  &  '0'  &  x"20";	
		tmp(246) := LDA  &  R0  &  '1'  &  x"61";	
		tmp(247) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(248) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(249) := LDA  &  R2  &  '1'  &  x"40";	
		tmp(250) := JEQ  &  R0  &  '0'  &  x"f4";	
		tmp(251) := STA  &  R2  &  '0'  &  x"0f";	
		tmp(252) := STA  &  R2  &  '1'  &  x"25";	
		tmp(253) := STA  &  R0  &  '1'  &  x"fe";	
		tmp(254) := LDA  &  R3  &  '0'  &  x"07";	
		tmp(256) := LDA  &  R0  &  '0'  &  x"0e";	
		tmp(257) := LDA  &  R1  &  '0'  &  x"0f";	
		tmp(258) := LDA  &  R2  &  '0'  &  x"07";	
		tmp(259) := ADDI  &  R3  &  '0'  &  x"0a";	
		tmp(261) := CEQ  &  R1  &  '0'  &  x"07";	
		tmp(262) := JEQ  &  R0  &  '1'  &  x"08";	
		tmp(263) := JMP  &  R0  &  '1'  &  x"03";	
		tmp(264) := SOMA  &  R3  &  '0'  &  x"0e";	
		tmp(265) := CLT  &  R3  &  '0'  &  x"13";	
		tmp(266) := JLT  &  R0  &  '1'  &  x"25";	
		tmp(267) := CEQ  &  R3  &  '0'  &  x"13";	
		tmp(268) := JEQ  &  R0  &  '1'  &  x"10";	
		tmp(269) := LDA  &  R0  &  '0'  &  x"08";	
		tmp(271) := JMP  &  R0  &  '0'  &  x"c2";	
		tmp(272) := LDA  &  R0  &  '0'  &  x"08";	
		tmp(274) := LDA  &  R0  &  '0'  &  x"07";	
		tmp(275) := STA  &  R0  &  '0'  &  x"0e";	
		tmp(276) := STA  &  R0  &  '0'  &  x"0f";	
		tmp(277) := LDA  &  R0  &  '0'  &  x"0a";	
		tmp(278) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(279) := JEQ  &  R0  &  '1'  &  x"19";	
		tmp(280) := JMP  &  R0  &  '0'  &  x"c2";	
		tmp(281) := LDA  &  R0  &  '0'  &  x"0b";	
		tmp(282) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(283) := JEQ  &  R0  &  '1'  &  x"1d";	
		tmp(284) := JMP  &  R0  &  '0'  &  x"cc";	
		tmp(285) := LDA  &  R0  &  '0'  &  x"0c";	
		tmp(286) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(287) := JEQ  &  R0  &  '1'  &  x"21";	
		tmp(288) := JMP  &  R0  &  '0'  &  x"d6";	
		tmp(289) := LDA  &  R0  &  '0'  &  x"0d";	
		tmp(290) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(291) := JEQ  &  R0  &  '1'  &  x"25";	
		tmp(292) := JMP  &  R0  &  '0'  &  x"e0";	
		tmp(293) := LDA  &  R0  &  '0'  &  x"07";	
		tmp(295) := RET  &  R0  &  '0'  &  x"00";	
		tmp(296) := STA  &  R0  &  '1'  &  x"fd";	
		tmp(297) := LDA  &  R0  &  '0'  &  x"07";	
		tmp(301) := LDA  &  R2  &  '0'  &  x"10";	
		tmp(308) := RET  &  R0  &  '0'  &  x"00";	
		tmp(309) := STA  &  R0  &  '1'  &  x"fc";	
		tmp(310) := LDA  &  R1  &  '0'  &  x"08";	
		tmp(312) := LDA  &  R0  &  '1'  &  x"63";	
		tmp(313) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(314) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(315) := LDA  &  R2  &  '1'  &  x"40";	
		tmp(316) := JEQ  &  R0  &  '1'  &  x"36";	
		tmp(317) := STA  &  R2  &  '0'  &  x"00";	
		tmp(318) := STA  &  R2  &  '1'  &  x"20";	
		tmp(319) := STA  &  R0  &  '1'  &  x"fc";	
		tmp(320) := LDI  &  R1  &  '0'  &  x"02";	
		tmp(322) := LDA  &  R0  &  '1'  &  x"63";	
		tmp(323) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(324) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(325) := LDA  &  R2  &  '1'  &  x"40";	
		tmp(326) := JEQ  &  R0  &  '1'  &  x"40";	
		tmp(327) := STA  &  R2  &  '0'  &  x"01";	
		tmp(328) := STA  &  R2  &  '1'  &  x"21";	
		tmp(329) := STA  &  R0  &  '1'  &  x"fc";	
		tmp(330) := LDI  &  R1  &  '0'  &  x"04";	
		tmp(332) := LDA  &  R0  &  '1'  &  x"63";	
		tmp(333) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(334) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(335) := LDA  &  R2  &  '1'  &  x"40";	
		tmp(336) := JEQ  &  R0  &  '1'  &  x"4a";	
		tmp(337) := STA  &  R2  &  '0'  &  x"02";	
		tmp(338) := STA  &  R2  &  '1'  &  x"22";	
		tmp(339) := STA  &  R0  &  '1'  &  x"fc";	
		tmp(340) := LDI  &  R1  &  '0'  &  x"08";	
		tmp(342) := LDA  &  R0  &  '1'  &  x"63";	
		tmp(343) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(344) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(345) := LDA  &  R2  &  '1'  &  x"40";	
		tmp(346) := JEQ  &  R0  &  '1'  &  x"54";	
		tmp(347) := STA  &  R2  &  '0'  &  x"03";	
		tmp(348) := STA  &  R2  &  '1'  &  x"23";	
		tmp(349) := STA  &  R0  &  '1'  &  x"fc";	
		tmp(350) := LDI  &  R1  &  '0'  &  x"10";	
		tmp(352) := LDA  &  R0  &  '1'  &  x"63";	
		tmp(353) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(354) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(355) := LDA  &  R2  &  '1'  &  x"40";	
		tmp(356) := JEQ  &  R0  &  '1'  &  x"5e";	
		tmp(357) := STA  &  R2  &  '0'  &  x"04";	
		tmp(358) := STA  &  R2  &  '1'  &  x"24";	
		tmp(359) := STA  &  R0  &  '1'  &  x"fc";	
		tmp(360) := LDI  &  R1  &  '0'  &  x"20";	
		tmp(362) := LDA  &  R0  &  '1'  &  x"63";	
		tmp(363) := ANDI  &  R0  &  '0'  &  x"01";	
		tmp(364) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(365) := LDA  &  R2  &  '1'  &  x"40";	
		tmp(366) := JEQ  &  R0  &  '1'  &  x"68";	
		tmp(367) := STA  &  R2  &  '0'  &  x"05";	
		tmp(368) := STA  &  R2  &  '1'  &  x"25";	
		tmp(369) := STA  &  R0  &  '1'  &  x"fc";	
		tmp(370) := LDA  &  R3  &  '0'  &  x"07";	
		tmp(372) := LDA  &  R0  &  '0'  &  x"04";	
		tmp(373) := LDA  &  R1  &  '0'  &  x"05";	
		tmp(374) := LDA  &  R2  &  '0'  &  x"07";	
		tmp(375) := ADDI  &  R3  &  '0'  &  x"0a";	
		tmp(377) := CEQ  &  R1  &  '0'  &  x"07";	
		tmp(378) := JEQ  &  R0  &  '1'  &  x"7c";	
		tmp(379) := JMP  &  R0  &  '1'  &  x"77";	
		tmp(380) := SOMA  &  R3  &  '0'  &  x"04";	
		tmp(381) := CLT  &  R3  &  '0'  &  x"13";	
		tmp(382) := JLT  &  R0  &  '1'  &  x"99";	
		tmp(383) := CEQ  &  R3  &  '0'  &  x"13";	
		tmp(384) := JEQ  &  R0  &  '1'  &  x"84";	
		tmp(385) := LDA  &  R0  &  '0'  &  x"08";	
		tmp(387) := JMP  &  R0  &  '1'  &  x"36";	
		tmp(388) := LDA  &  R0  &  '0'  &  x"08";	
		tmp(390) := LDA  &  R0  &  '0'  &  x"07";	
		tmp(391) := STA  &  R0  &  '0'  &  x"04";	
		tmp(392) := STA  &  R0  &  '0'  &  x"05";	
		tmp(393) := LDA  &  R0  &  '0'  &  x"00";	
		tmp(394) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(395) := JEQ  &  R0  &  '1'  &  x"8d";	
		tmp(396) := JMP  &  R0  &  '1'  &  x"36";	
		tmp(397) := LDA  &  R0  &  '0'  &  x"01";	
		tmp(398) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(399) := JEQ  &  R0  &  '1'  &  x"91";	
		tmp(400) := JMP  &  R0  &  '1'  &  x"40";	
		tmp(401) := LDA  &  R0  &  '0'  &  x"02";	
		tmp(402) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(403) := JEQ  &  R0  &  '1'  &  x"95";	
		tmp(404) := JMP  &  R0  &  '1'  &  x"4a";	
		tmp(405) := LDA  &  R0  &  '0'  &  x"03";	
		tmp(406) := CEQ  &  R0  &  '0'  &  x"07";	
		tmp(407) := JEQ  &  R0  &  '1'  &  x"99";	
		tmp(408) := JMP  &  R0  &  '1'  &  x"54";	
		tmp(409) := LDA  &  R0  &  '0'  &  x"07";	
		tmp(411) := RET  &  R0  &  '0'  &  x"00";	

		  return tmp;
		  
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;